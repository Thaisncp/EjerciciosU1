--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity promedio1 is
	Port ( A, B : in STD_LOGIC_VECTOR ( 2 downto 0); 
			C : out STD_LOGIC_VECTOR (2 downto 0)); 
end promedio1;


