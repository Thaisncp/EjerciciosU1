--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiplexor2 is
	Port ( E0, E1, E2, E3 : in  STD_LOGIC_VECTOR(0 to 3);
          S0, S1 : in  STD_LOGIC_VECTOR(0 to 3);
          F : out  STD_LOGIC);
end multiplexor2;


