--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidadB is
    Port ( P0, P1, P2 : in  STD_LOGIC;
           A0, A1 : out  STD_LOGIC);
end entidadB;

