--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity promedio2 is
	Port ( A, B : in STD_LOGIC_VECTOR ( 0 to 3 );
			C : out STD_LOGIC_VECTOR (0 to 3 )) ;
end promedio2;
