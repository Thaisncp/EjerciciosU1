--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidadA is
    Port ( A, B : in  STD_LOGIC;
           C : out  STD_LOGIC);
end entidadA;

