--Thais Cartuche
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiplexor is
	Port ( E0 , El, E2 , E3 : in STD_LOGIC; 
			S0 , Sl : in STD_LOGIC ;
			F : out STD_LOGIC);
end multiplexor;

